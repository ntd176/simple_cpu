`timescale 1ns / 1ns

module cpu_tb;
    reg        clk_tb;
    reg        resetn_tb;
    reg        run_tb;
    reg [15:0] din_tb;
    wire       done_tb;

    cpu dut (
        .clk(clk_tb),
        .resetn(resetn_tb),
        .run(run_tb),
        .din(din_tb),
        .done(done_tb)
    );

    initial begin
        clk_tb = 0;
        forever #10 clk_tb = ~clk_tb;
    end

    localparam MV  = 3'b000;
    localparam MVI = 3'b001;
    localparam ADD = 3'b010;
    localparam SUB = 3'b011;

    initial begin
        run_tb    = 1'b1;
        din_tb    = 16'hXXXX;
        resetn_tb = 1'b1;
        #40;
		run_tb = 1'b0; // off system
        #60;
		run_tb = 1'b1;
		resetn_tb = 1'b0; // reset system
        #20;
		resetn_tb = 1'b1;
		
        //---MVI---//
		//--mvi, r0, 000Ah--//
        din_tb = {7'b0, MVI, 3'd0, 3'd0}; // State 0 --> instruction fetch
        #20;
        din_tb = 16'h000A;                // State 1 --> data fetch
        #20;
		//-------------------------------
		//--mvi, r1, 0008h--//
        din_tb = {7'b0, MVI, 3'd1, 3'd0};
        #20;
        din_tb = 16'h0008;
        #20;
		//-------------------------------
		//--mvi, r2, 0006h--//
        din_tb = {7'b0, MVI, 3'd2, 3'd0};
        #20;
        din_tb = 16'h0006;
        #20;
		//-------------------------------
		//--mvi, r3, 0002h--//
        din_tb = {7'b0, MVI, 3'd3, 3'd0};
        #20;
        din_tb = 16'h0002;
        #20;
		//-------------------------------
		//--mvi, r4, FFFFh--//
        din_tb = {7'b0, MVI, 3'd4, 3'd0};
        #20;
        din_tb = 16'hFFFF;
        #20;
		//-------------------------------
		//--mvi, r5, EEEEh--//
        din_tb = {7'b0, MVI, 3'd5, 3'd0};
        #20;
        din_tb = 16'hEEEE;
        #20;
		//-------------------------------
		//--mvi, r6, CCCCh--//
        din_tb = {7'b0, MVI, 3'd6, 3'd0};
        #20;
        din_tb = 16'hCCCC;
        #20;
		//-------------------------------
		//--mvi, r7, DDDDh--//
        din_tb = {7'b0, MVI, 3'd7, 3'd0};
        #20;
        din_tb = 16'hDDDD;
        #20;
		//=================================
		//---MV---//
		//--mv, r7, r0--//
        din_tb = {7'b0, MV, 3'd7, 3'd0};
        #20;
        din_tb = 16'h000A;
        #20;
		//-------------------------------
		//--mv, r6, r1--//
        din_tb = {7'b0, MV, 3'd6, 3'd1};
        #20;
        din_tb = 16'h0008;
        #20;
		//-------------------------------
		//--mv, r5, r2--//
        din_tb = {7'b0, MV, 3'd5, 3'd2};
        #20;
        din_tb = 16'h0006;
        #20;
		//-------------------------------
		//--mv, r4, r3--//
        din_tb = {7'b0, MV, 3'd4, 3'd3};
        #20;
        din_tb = 16'h0002;
        #20;
		//-------------------------------
		//--mv, r3, r7--//
        din_tb = {7'b0, MV, 3'd3, 3'd7};
        #20;
        din_tb = 16'h000A;
        #20;
		//-------------------------------
		//--mv, r2, r6 --//
        din_tb = {7'b0, MV, 3'd2, 3'd6};
        #20;
        din_tb = 16'h0008;
        #20;
		//-------------------------------
		//--mv, r1, r5--//
        din_tb = {7'b0, MV, 3'd1, 3'd5};
        #20;
        din_tb = 16'h0006;
        #20;
		//-------------------------------
		//--mv, r0, r4--//
        din_tb = {7'b0, MV, 3'd0, 3'd4};
        #20;
        din_tb = 16'h0002;
        #20;
		//=================================
		//---ADD---//
		//--add, r0, r1--//
        din_tb = {7'b0, ADD, 3'd0, 3'd1};	// fetch
        #20;
        // load A
        #20;
		// execute
		#20;
		// writeback
		#20;	// result r0 = 0008h
		//-------------------------------
		//--add, r1, r2--//
        din_tb = {7'b0, ADD, 3'd1, 3'd2};
        #20;
        #20;
		#20;
		#20;	// result r1 = 000Eh
		//-------------------------------
		//--add, r2, r3--//
        din_tb = {7'b0, ADD, 3'd2, 3'd3};
        #20;
        #20;
		#20;
		#20;	// result r2 = 0012h
		//-------------------------------
		//--add, r3, r4--//
        din_tb = {7'b0, ADD, 3'd3, 3'd4};
        #20;
        #20;
		#20;
		#20;	// result r3 = 000Ch
		//-------------------------------
		//--add, r4, r5--//
        din_tb = {7'b0, ADD, 3'd4, 3'd5};
        #20;
        #20;
		#20;
		#20;	// result r4 = 0008h
		//-------------------------------
		//--add, r5, r6--//
        din_tb = {7'b0, ADD, 3'd5, 3'd6};
        #20;
        #20;
		#20;
		#20;	// result r5 = 000Eh
		//-------------------------------
		//--add, r6, r7--//
        din_tb = {7'b0, ADD, 3'd6, 3'd7};
        #20;
        #20;
		#20;
		#20;	// result r6 = 0012h
		//-------------------------------
		//--add, r7, r1--//
        din_tb = {7'b0, ADD, 3'd7, 3'd1};
        #20;
        #20;
		#20;
		#20;	// result r7 = 0012h
		//-------------------------------
		//=================================
		//---SUB---//
		//--sub, r7, r6--//
        din_tb = {7'b0, SUB, 3'd7, 3'd6};
        #20;
        #20;
		#20;
		#20;	// result r7 = 0000h
		//-------------------------------
		//--sub, r6, r5--//
        din_tb = {7'b0, SUB, 3'd6, 3'd5};
        #20;
        #20;
		#20;
		#20;	// result r6 = 0004h
		//-------------------------------
		//--sub, r5, r4--//
        din_tb = {7'b0, SUB, 3'd5, 3'd4};
        #20;
        #20;
		#20;
		#20;	// result r5 = 0006h
		//-------------------------------
		//--sub, r3, r4--//
        din_tb = {7'b0, SUB, 3'd3, 3'd4};
        #20;
        #20;
		#20;
		#20;	// result r3 = 0004h
		//-------------------------------
		//--sub, r4, r3--//
        din_tb = {7'b0, SUB, 3'd4, 3'd3};
        #20;
        #20;
		#20;
		#20;	// result r4 = 0004h
		//-------------------------------
		//--sub, r2, r3--//
        din_tb = {7'b0, SUB, 3'd2, 3'd3};
        #20;
        #20;
		#20;
		#20;	// result r2 = 0006h
		//-------------------------------
		//--sub, r1, r0--//
        din_tb = {7'b0, SUB, 3'd1, 3'd0};
        #20;
        #20;
		#20;
		#20;	// result r1 = 0006h
		//-------------------------------
		//--sub, r0, r1--//
        din_tb = {7'b0, SUB, 3'd0, 3'd1};
        #20;
        #20;
		#20;
		#20;	// result r0 = 0002h
		//-------------------------------
        $finish;
    end
	
endmodule